`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:24:02 11/15/2017 
// Design Name: 
// Module Name:    huffman 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module huffman(
						A11, A12, A13, A14, A15, A16, A17, A18,
						A21, A22, A23, A24, A25, A26, A27, A28,
						A31, A32, A33, A34, A35, A36, A37, A38,
						A41, A42, A43, A44, A45, A46, A47, A48,
						A51, A52, A53, A54, A55, A56, A57, A58,
						A61, A62, A63, A64, A65, A66, A67, A68,
						A71, A72, A73, A74, A75, A76, A77, A78,
						A81, A82, A83, A84, A85, A86, A87, A88,
						
						B11, B12, B13, B14, B15, B16, B17, B18,
						B21, B22, B23, B24, B25, B26, B27, B28,
						B31, B32, B33, B34, B35, B36, B37, B38,
						B41, B42, B43, B44, B45, B46, B47, B48,
						B51, B52, B53, B54, B55, B56, B57, B58,
						B61, B62, B63, B64, B65, B66, B67, B68,
						B71, B72, B73, B74, B75, B76, B77, B78,
						B81, B82, B83, B84, B85, B86, B87, B88,
    );

input [31:0] A11, A12, A13, A14, A15, A16, A17, A18,
					 A21, A22, A23, A24, A25, A26, A27, A28,
					 A31, A32, A33, A34, A35, A36, A37, A38,
					 A41, A42, A43, A44, A45, A46, A47, A48,
					 A51, A52, A53, A54, A55, A56, A57, A58,
					 A61, A62, A63, A64, A65, A66, A67, A68,
					 A71, A72, A73, A74, A75, A76, A77, A78,
					 A81, A82, A83, A84, A85, A86, A87, A88;
					 
	output [15:0] B11, B12, B13, B14, B15, B16, B17, B18,
					 B21, B22, B23, B24, B25, B26, B27, B28,
					 B31, B32, B33, B34, B35, B36, B37, B38,
					 B41, B42, B43, B44, B45, B46, B47, B48,
					 B51, B52, B53, B54, B55, B56, B57, B58,
					 B61, B62, B63, B64, B65, B66, B67, B68,
					 B71, B72, B73, B74, B75, B76, B77, B78,
					 B81, B82, B83, B84, B85, B86, B87, B88;
					 
					 assign B11 = (A11[31:16] == 0)?0:
					             (A11[31:16] == 16'b0000_0000_0000_0001)?16'b0000_0000_0000_0001:
									 (A11[31:16] == 16'b0000_0000_0000_0010)?16'b0000_0000_0000_1000:
									 (A11[31:16] == 16'b0000_0000_0000_0011)?16'b0000_0000_0000_1001:
									 (A11[31:16] == 16'b0000_0000_0000_0100)?16'b0000_0000_0000_1010:
									 (A11[31:16] == 16'b0000_0000_0000_0101)?16'b0000_0000_0000_1011:
									 (A11[31:16] == 16'b0000_0000_0000_0110)?16'b0000_0000_0000_1100:
									 (A11[31:16] == 16'b0000_0000_0000_0111)?16'b0000_0000_0000_1101:
									 (A11[31:16] == 16'b0000_0000_0000_1000)?16'b0000_0000_0001_1100:
									 (A11[31:16] == 16'b0000_0000_0000_1001)?16'b0000_0000_0011_1010:
									 (A11[31:16] == 16'b0000_0000_0000_1010)?16'b0000_0000_0011_1011:
									 (A11[31:16] == 16'b0000_0000_0000_1011)?16'b0000_0000_0011_1100:
									 (A11[31:16] == 16'b0000_0000_0000_1100)?16'b0000_0000_0111_1010:
									 (A11[31:16] == 16'b0000_0000_0000_1101)?16'b0000_0000_0111_1011:
									 (A11[31:16] == 16'b0000_0000_0000_1110)?16'b0000_0000_1111_1000:
									 (A11[31:16] == 16'b0000_0000_0000_1111)?16'b0000_0000_1111_1001:
									 (A11[31:16] == 16'b0000_0000_0001_0000)?16'b0000_0000_1111_1010:
									 (A11[31:16] == 16'b0000_0000_0001_0001)?16'b0000_0000_1111_1011:
									 (A11[31:16] == 16'b0000_0000_0001_0010)?16'b0000_0000_1111_1100:
									 (A11[31:16] == 16'b0000_0000_0001_0011)?16'b0000_0001_1111_1010:
									 (A11[31:16] == 16'b0000_0000_0001_0100)?16'b0000_0001_1111_1011:
									 (A11[31:16] == 16'b0000_0000_0001_0101)?16'b0000_0001_1111_1100:
									 (A11[31:16] == 16'b0000_0000_0001_0110)?16'b0000_0011_1111_1010:
									 (A11[31:16] == 16'b0000_0000_0001_0111)?16'b0000_0011_1111_1011:
									 (A11[31:16] == 16'b0000_0000_0001_1000)?16'b0000_0011_1111_1100:
									 (A11[31:16] == 16'b0000_0000_0001_1001)?16'b0000_0011_1111_1101:
									 (A11[31:16] == 16'b0000_0000_0001_1010)?16'b0000_0011_1111_1110:
									 (A11[31:16] == 16'b0000_0000_0001_1011)?16'b0000_1111_1111_1100:
									 (A11[31:16] == 16'b0000_0000_0001_1100)?16'b0000_1111_1111_1101:
									 (A11[31:16] == 16'b0000_0000_0001_1101)?16'b0000_1111_1111_1110:
									 (A11[31:16] == 16'b0000_0000_0001_1110)?16'b0001_1111_1111_1110:
									 (A11[31:16] == 16'b0000_0000_0001_1111)?16'b0001_1111_1111_1111:16'b1111_1111_1111_1111;
endmodule
